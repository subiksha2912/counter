module counter_tb.v;
  
